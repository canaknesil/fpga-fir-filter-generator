
library IEEE; 
use IEEE.STD_LOGIC_1164.ALL; 

entity threesamplefilter is 
	Port ( input : in  STD_LOGIC_VECTOR (7 downto 0); 
		clock : in  STD_LOGIC; 
		output : out  STD_LOGIC_VECTOR (7 downto 0)); 
end threesamplefilter; 

architecture Behavioral of threesamplefilter is 

component module1 is 
	Port ( input : in  STD_LOGIC_VECTOR (7 downto 0); 
		term : in  STD_LOGIC_VECTOR (7 downto 0); 
		hardcoded : in std_logic_vector (7 downto 0); 
		output : out  STD_LOGIC_VECTOR (7 downto 0)); 
end component; 

component module2 is 
	Port ( input : in  STD_LOGIC_VECTOR (7 downto 0); 
		term : in  STD_LOGIC_VECTOR (7 downto 0); 
		clock : in  STD_LOGIC; 
		hardcoded : in std_logic_vector (7 downto 0); 
		output : out  STD_LOGIC_VECTOR (7 downto 0); 
		fout : out  STD_LOGIC_VECTOR (7 downto 0)); 
end component; 

component module3 is 
	Port ( input : in  STD_LOGIC_VECTOR (7 downto 0); 
		clock : in  STD_LOGIC; 
		hardcoded : in std_logic_vector (7 downto 0); 
		output : out  STD_LOGIC_VECTOR (7 downto 0)); 
end component; 

signal hardcoded_0: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_1: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_2: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_3: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_4: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_5: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_6: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_7: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_8: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_9: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_10: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_11: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_12: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_13: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_14: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_15: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_16: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_17: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_18: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_19: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_20: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_21: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_22: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_23: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_24: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_25: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_26: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_27: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_28: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_29: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_30: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_31: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_32: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_33: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_34: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_35: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_36: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_37: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_38: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_39: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_40: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_41: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_42: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_43: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_44: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_45: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_46: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_47: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_48: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_49: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_50: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_51: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_52: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_53: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_54: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_55: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_56: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_57: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_58: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_59: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_60: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_61: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_62: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_63: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_64: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_65: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_66: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_67: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_68: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_69: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_70: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_71: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_72: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_73: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_74: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_75: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_76: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_77: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_78: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_79: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_80: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_81: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_82: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_83: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_84: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_85: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_86: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_87: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_88: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_89: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_90: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_91: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_92: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_93: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_94: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_95: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_96: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_97: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_98: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_99: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_100: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_101: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_102: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_103: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_104: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_105: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_106: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_107: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_108: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_109: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_110: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_111: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_112: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_113: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_114: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_115: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_116: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_117: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_118: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_119: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_120: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_121: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_122: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_123: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_124: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_125: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_126: std_logic_vector(7 downto 0) := "00000001"; 
signal hardcoded_127: std_logic_vector(7 downto 0) := "00000001"; 

signal module1_term: std_logic_vector(7 downto 0); 

signal module2_1_todown, module2_1_fromdown : std_logic_vector(7 downto 0); 
signal module2_2_todown, module2_2_fromdown : std_logic_vector(7 downto 0); 
signal module2_3_todown, module2_3_fromdown : std_logic_vector(7 downto 0); 
signal module2_4_todown, module2_4_fromdown : std_logic_vector(7 downto 0); 
signal module2_5_todown, module2_5_fromdown : std_logic_vector(7 downto 0); 
signal module2_6_todown, module2_6_fromdown : std_logic_vector(7 downto 0); 
signal module2_7_todown, module2_7_fromdown : std_logic_vector(7 downto 0); 
signal module2_8_todown, module2_8_fromdown : std_logic_vector(7 downto 0); 
signal module2_9_todown, module2_9_fromdown : std_logic_vector(7 downto 0); 
signal module2_10_todown, module2_10_fromdown : std_logic_vector(7 downto 0); 
signal module2_11_todown, module2_11_fromdown : std_logic_vector(7 downto 0); 
signal module2_12_todown, module2_12_fromdown : std_logic_vector(7 downto 0); 
signal module2_13_todown, module2_13_fromdown : std_logic_vector(7 downto 0); 
signal module2_14_todown, module2_14_fromdown : std_logic_vector(7 downto 0); 
signal module2_15_todown, module2_15_fromdown : std_logic_vector(7 downto 0); 
signal module2_16_todown, module2_16_fromdown : std_logic_vector(7 downto 0); 
signal module2_17_todown, module2_17_fromdown : std_logic_vector(7 downto 0); 
signal module2_18_todown, module2_18_fromdown : std_logic_vector(7 downto 0); 
signal module2_19_todown, module2_19_fromdown : std_logic_vector(7 downto 0); 
signal module2_20_todown, module2_20_fromdown : std_logic_vector(7 downto 0); 
signal module2_21_todown, module2_21_fromdown : std_logic_vector(7 downto 0); 
signal module2_22_todown, module2_22_fromdown : std_logic_vector(7 downto 0); 
signal module2_23_todown, module2_23_fromdown : std_logic_vector(7 downto 0); 
signal module2_24_todown, module2_24_fromdown : std_logic_vector(7 downto 0); 
signal module2_25_todown, module2_25_fromdown : std_logic_vector(7 downto 0); 
signal module2_26_todown, module2_26_fromdown : std_logic_vector(7 downto 0); 
signal module2_27_todown, module2_27_fromdown : std_logic_vector(7 downto 0); 
signal module2_28_todown, module2_28_fromdown : std_logic_vector(7 downto 0); 
signal module2_29_todown, module2_29_fromdown : std_logic_vector(7 downto 0); 
signal module2_30_todown, module2_30_fromdown : std_logic_vector(7 downto 0); 
signal module2_31_todown, module2_31_fromdown : std_logic_vector(7 downto 0); 
signal module2_32_todown, module2_32_fromdown : std_logic_vector(7 downto 0); 
signal module2_33_todown, module2_33_fromdown : std_logic_vector(7 downto 0); 
signal module2_34_todown, module2_34_fromdown : std_logic_vector(7 downto 0); 
signal module2_35_todown, module2_35_fromdown : std_logic_vector(7 downto 0); 
signal module2_36_todown, module2_36_fromdown : std_logic_vector(7 downto 0); 
signal module2_37_todown, module2_37_fromdown : std_logic_vector(7 downto 0); 
signal module2_38_todown, module2_38_fromdown : std_logic_vector(7 downto 0); 
signal module2_39_todown, module2_39_fromdown : std_logic_vector(7 downto 0); 
signal module2_40_todown, module2_40_fromdown : std_logic_vector(7 downto 0); 
signal module2_41_todown, module2_41_fromdown : std_logic_vector(7 downto 0); 
signal module2_42_todown, module2_42_fromdown : std_logic_vector(7 downto 0); 
signal module2_43_todown, module2_43_fromdown : std_logic_vector(7 downto 0); 
signal module2_44_todown, module2_44_fromdown : std_logic_vector(7 downto 0); 
signal module2_45_todown, module2_45_fromdown : std_logic_vector(7 downto 0); 
signal module2_46_todown, module2_46_fromdown : std_logic_vector(7 downto 0); 
signal module2_47_todown, module2_47_fromdown : std_logic_vector(7 downto 0); 
signal module2_48_todown, module2_48_fromdown : std_logic_vector(7 downto 0); 
signal module2_49_todown, module2_49_fromdown : std_logic_vector(7 downto 0); 
signal module2_50_todown, module2_50_fromdown : std_logic_vector(7 downto 0); 
signal module2_51_todown, module2_51_fromdown : std_logic_vector(7 downto 0); 
signal module2_52_todown, module2_52_fromdown : std_logic_vector(7 downto 0); 
signal module2_53_todown, module2_53_fromdown : std_logic_vector(7 downto 0); 
signal module2_54_todown, module2_54_fromdown : std_logic_vector(7 downto 0); 
signal module2_55_todown, module2_55_fromdown : std_logic_vector(7 downto 0); 
signal module2_56_todown, module2_56_fromdown : std_logic_vector(7 downto 0); 
signal module2_57_todown, module2_57_fromdown : std_logic_vector(7 downto 0); 
signal module2_58_todown, module2_58_fromdown : std_logic_vector(7 downto 0); 
signal module2_59_todown, module2_59_fromdown : std_logic_vector(7 downto 0); 
signal module2_60_todown, module2_60_fromdown : std_logic_vector(7 downto 0); 
signal module2_61_todown, module2_61_fromdown : std_logic_vector(7 downto 0); 
signal module2_62_todown, module2_62_fromdown : std_logic_vector(7 downto 0); 
signal module2_63_todown, module2_63_fromdown : std_logic_vector(7 downto 0); 
signal module2_64_todown, module2_64_fromdown : std_logic_vector(7 downto 0); 
signal module2_65_todown, module2_65_fromdown : std_logic_vector(7 downto 0); 
signal module2_66_todown, module2_66_fromdown : std_logic_vector(7 downto 0); 
signal module2_67_todown, module2_67_fromdown : std_logic_vector(7 downto 0); 
signal module2_68_todown, module2_68_fromdown : std_logic_vector(7 downto 0); 
signal module2_69_todown, module2_69_fromdown : std_logic_vector(7 downto 0); 
signal module2_70_todown, module2_70_fromdown : std_logic_vector(7 downto 0); 
signal module2_71_todown, module2_71_fromdown : std_logic_vector(7 downto 0); 
signal module2_72_todown, module2_72_fromdown : std_logic_vector(7 downto 0); 
signal module2_73_todown, module2_73_fromdown : std_logic_vector(7 downto 0); 
signal module2_74_todown, module2_74_fromdown : std_logic_vector(7 downto 0); 
signal module2_75_todown, module2_75_fromdown : std_logic_vector(7 downto 0); 
signal module2_76_todown, module2_76_fromdown : std_logic_vector(7 downto 0); 
signal module2_77_todown, module2_77_fromdown : std_logic_vector(7 downto 0); 
signal module2_78_todown, module2_78_fromdown : std_logic_vector(7 downto 0); 
signal module2_79_todown, module2_79_fromdown : std_logic_vector(7 downto 0); 
signal module2_80_todown, module2_80_fromdown : std_logic_vector(7 downto 0); 
signal module2_81_todown, module2_81_fromdown : std_logic_vector(7 downto 0); 
signal module2_82_todown, module2_82_fromdown : std_logic_vector(7 downto 0); 
signal module2_83_todown, module2_83_fromdown : std_logic_vector(7 downto 0); 
signal module2_84_todown, module2_84_fromdown : std_logic_vector(7 downto 0); 
signal module2_85_todown, module2_85_fromdown : std_logic_vector(7 downto 0); 
signal module2_86_todown, module2_86_fromdown : std_logic_vector(7 downto 0); 
signal module2_87_todown, module2_87_fromdown : std_logic_vector(7 downto 0); 
signal module2_88_todown, module2_88_fromdown : std_logic_vector(7 downto 0); 
signal module2_89_todown, module2_89_fromdown : std_logic_vector(7 downto 0); 
signal module2_90_todown, module2_90_fromdown : std_logic_vector(7 downto 0); 
signal module2_91_todown, module2_91_fromdown : std_logic_vector(7 downto 0); 
signal module2_92_todown, module2_92_fromdown : std_logic_vector(7 downto 0); 
signal module2_93_todown, module2_93_fromdown : std_logic_vector(7 downto 0); 
signal module2_94_todown, module2_94_fromdown : std_logic_vector(7 downto 0); 
signal module2_95_todown, module2_95_fromdown : std_logic_vector(7 downto 0); 
signal module2_96_todown, module2_96_fromdown : std_logic_vector(7 downto 0); 
signal module2_97_todown, module2_97_fromdown : std_logic_vector(7 downto 0); 
signal module2_98_todown, module2_98_fromdown : std_logic_vector(7 downto 0); 
signal module2_99_todown, module2_99_fromdown : std_logic_vector(7 downto 0); 
signal module2_100_todown, module2_100_fromdown : std_logic_vector(7 downto 0); 
signal module2_101_todown, module2_101_fromdown : std_logic_vector(7 downto 0); 
signal module2_102_todown, module2_102_fromdown : std_logic_vector(7 downto 0); 
signal module2_103_todown, module2_103_fromdown : std_logic_vector(7 downto 0); 
signal module2_104_todown, module2_104_fromdown : std_logic_vector(7 downto 0); 
signal module2_105_todown, module2_105_fromdown : std_logic_vector(7 downto 0); 
signal module2_106_todown, module2_106_fromdown : std_logic_vector(7 downto 0); 
signal module2_107_todown, module2_107_fromdown : std_logic_vector(7 downto 0); 
signal module2_108_todown, module2_108_fromdown : std_logic_vector(7 downto 0); 
signal module2_109_todown, module2_109_fromdown : std_logic_vector(7 downto 0); 
signal module2_110_todown, module2_110_fromdown : std_logic_vector(7 downto 0); 
signal module2_111_todown, module2_111_fromdown : std_logic_vector(7 downto 0); 
signal module2_112_todown, module2_112_fromdown : std_logic_vector(7 downto 0); 
signal module2_113_todown, module2_113_fromdown : std_logic_vector(7 downto 0); 
signal module2_114_todown, module2_114_fromdown : std_logic_vector(7 downto 0); 
signal module2_115_todown, module2_115_fromdown : std_logic_vector(7 downto 0); 
signal module2_116_todown, module2_116_fromdown : std_logic_vector(7 downto 0); 
signal module2_117_todown, module2_117_fromdown : std_logic_vector(7 downto 0); 
signal module2_118_todown, module2_118_fromdown : std_logic_vector(7 downto 0); 
signal module2_119_todown, module2_119_fromdown : std_logic_vector(7 downto 0); 
signal module2_120_todown, module2_120_fromdown : std_logic_vector(7 downto 0); 
signal module2_121_todown, module2_121_fromdown : std_logic_vector(7 downto 0); 
signal module2_122_todown, module2_122_fromdown : std_logic_vector(7 downto 0); 
signal module2_123_todown, module2_123_fromdown : std_logic_vector(7 downto 0); 
signal module2_124_todown, module2_124_fromdown : std_logic_vector(7 downto 0); 
signal module2_125_todown, module2_125_fromdown : std_logic_vector(7 downto 0); 
signal module2_126_todown, module2_126_fromdown : std_logic_vector(7 downto 0); 

begin 

module1op: module1 PORT MAP(input, module1_term, hardcoded_0, output); 
module2op_1: module2 PORT MAP(input, module2_1_fromdown, clock, hardcoded_1, module1_term, module2_1_todown); 
module2op_2: module2 PORT MAP(module2_1_todown, module2_2_fromdown, clock, hardcoded_2, module2_1_fromdown, module2_2_todown); 
module2op_3: module2 PORT MAP(module2_2_todown, module2_3_fromdown, clock, hardcoded_3, module2_2_fromdown, module2_3_todown); 
module2op_4: module2 PORT MAP(module2_3_todown, module2_4_fromdown, clock, hardcoded_4, module2_3_fromdown, module2_4_todown); 
module2op_5: module2 PORT MAP(module2_4_todown, module2_5_fromdown, clock, hardcoded_5, module2_4_fromdown, module2_5_todown); 
module2op_6: module2 PORT MAP(module2_5_todown, module2_6_fromdown, clock, hardcoded_6, module2_5_fromdown, module2_6_todown); 
module2op_7: module2 PORT MAP(module2_6_todown, module2_7_fromdown, clock, hardcoded_7, module2_6_fromdown, module2_7_todown); 
module2op_8: module2 PORT MAP(module2_7_todown, module2_8_fromdown, clock, hardcoded_8, module2_7_fromdown, module2_8_todown); 
module2op_9: module2 PORT MAP(module2_8_todown, module2_9_fromdown, clock, hardcoded_9, module2_8_fromdown, module2_9_todown); 
module2op_10: module2 PORT MAP(module2_9_todown, module2_10_fromdown, clock, hardcoded_10, module2_9_fromdown, module2_10_todown); 
module2op_11: module2 PORT MAP(module2_10_todown, module2_11_fromdown, clock, hardcoded_11, module2_10_fromdown, module2_11_todown); 
module2op_12: module2 PORT MAP(module2_11_todown, module2_12_fromdown, clock, hardcoded_12, module2_11_fromdown, module2_12_todown); 
module2op_13: module2 PORT MAP(module2_12_todown, module2_13_fromdown, clock, hardcoded_13, module2_12_fromdown, module2_13_todown); 
module2op_14: module2 PORT MAP(module2_13_todown, module2_14_fromdown, clock, hardcoded_14, module2_13_fromdown, module2_14_todown); 
module2op_15: module2 PORT MAP(module2_14_todown, module2_15_fromdown, clock, hardcoded_15, module2_14_fromdown, module2_15_todown); 
module2op_16: module2 PORT MAP(module2_15_todown, module2_16_fromdown, clock, hardcoded_16, module2_15_fromdown, module2_16_todown); 
module2op_17: module2 PORT MAP(module2_16_todown, module2_17_fromdown, clock, hardcoded_17, module2_16_fromdown, module2_17_todown); 
module2op_18: module2 PORT MAP(module2_17_todown, module2_18_fromdown, clock, hardcoded_18, module2_17_fromdown, module2_18_todown); 
module2op_19: module2 PORT MAP(module2_18_todown, module2_19_fromdown, clock, hardcoded_19, module2_18_fromdown, module2_19_todown); 
module2op_20: module2 PORT MAP(module2_19_todown, module2_20_fromdown, clock, hardcoded_20, module2_19_fromdown, module2_20_todown); 
module2op_21: module2 PORT MAP(module2_20_todown, module2_21_fromdown, clock, hardcoded_21, module2_20_fromdown, module2_21_todown); 
module2op_22: module2 PORT MAP(module2_21_todown, module2_22_fromdown, clock, hardcoded_22, module2_21_fromdown, module2_22_todown); 
module2op_23: module2 PORT MAP(module2_22_todown, module2_23_fromdown, clock, hardcoded_23, module2_22_fromdown, module2_23_todown); 
module2op_24: module2 PORT MAP(module2_23_todown, module2_24_fromdown, clock, hardcoded_24, module2_23_fromdown, module2_24_todown); 
module2op_25: module2 PORT MAP(module2_24_todown, module2_25_fromdown, clock, hardcoded_25, module2_24_fromdown, module2_25_todown); 
module2op_26: module2 PORT MAP(module2_25_todown, module2_26_fromdown, clock, hardcoded_26, module2_25_fromdown, module2_26_todown); 
module2op_27: module2 PORT MAP(module2_26_todown, module2_27_fromdown, clock, hardcoded_27, module2_26_fromdown, module2_27_todown); 
module2op_28: module2 PORT MAP(module2_27_todown, module2_28_fromdown, clock, hardcoded_28, module2_27_fromdown, module2_28_todown); 
module2op_29: module2 PORT MAP(module2_28_todown, module2_29_fromdown, clock, hardcoded_29, module2_28_fromdown, module2_29_todown); 
module2op_30: module2 PORT MAP(module2_29_todown, module2_30_fromdown, clock, hardcoded_30, module2_29_fromdown, module2_30_todown); 
module2op_31: module2 PORT MAP(module2_30_todown, module2_31_fromdown, clock, hardcoded_31, module2_30_fromdown, module2_31_todown); 
module2op_32: module2 PORT MAP(module2_31_todown, module2_32_fromdown, clock, hardcoded_32, module2_31_fromdown, module2_32_todown); 
module2op_33: module2 PORT MAP(module2_32_todown, module2_33_fromdown, clock, hardcoded_33, module2_32_fromdown, module2_33_todown); 
module2op_34: module2 PORT MAP(module2_33_todown, module2_34_fromdown, clock, hardcoded_34, module2_33_fromdown, module2_34_todown); 
module2op_35: module2 PORT MAP(module2_34_todown, module2_35_fromdown, clock, hardcoded_35, module2_34_fromdown, module2_35_todown); 
module2op_36: module2 PORT MAP(module2_35_todown, module2_36_fromdown, clock, hardcoded_36, module2_35_fromdown, module2_36_todown); 
module2op_37: module2 PORT MAP(module2_36_todown, module2_37_fromdown, clock, hardcoded_37, module2_36_fromdown, module2_37_todown); 
module2op_38: module2 PORT MAP(module2_37_todown, module2_38_fromdown, clock, hardcoded_38, module2_37_fromdown, module2_38_todown); 
module2op_39: module2 PORT MAP(module2_38_todown, module2_39_fromdown, clock, hardcoded_39, module2_38_fromdown, module2_39_todown); 
module2op_40: module2 PORT MAP(module2_39_todown, module2_40_fromdown, clock, hardcoded_40, module2_39_fromdown, module2_40_todown); 
module2op_41: module2 PORT MAP(module2_40_todown, module2_41_fromdown, clock, hardcoded_41, module2_40_fromdown, module2_41_todown); 
module2op_42: module2 PORT MAP(module2_41_todown, module2_42_fromdown, clock, hardcoded_42, module2_41_fromdown, module2_42_todown); 
module2op_43: module2 PORT MAP(module2_42_todown, module2_43_fromdown, clock, hardcoded_43, module2_42_fromdown, module2_43_todown); 
module2op_44: module2 PORT MAP(module2_43_todown, module2_44_fromdown, clock, hardcoded_44, module2_43_fromdown, module2_44_todown); 
module2op_45: module2 PORT MAP(module2_44_todown, module2_45_fromdown, clock, hardcoded_45, module2_44_fromdown, module2_45_todown); 
module2op_46: module2 PORT MAP(module2_45_todown, module2_46_fromdown, clock, hardcoded_46, module2_45_fromdown, module2_46_todown); 
module2op_47: module2 PORT MAP(module2_46_todown, module2_47_fromdown, clock, hardcoded_47, module2_46_fromdown, module2_47_todown); 
module2op_48: module2 PORT MAP(module2_47_todown, module2_48_fromdown, clock, hardcoded_48, module2_47_fromdown, module2_48_todown); 
module2op_49: module2 PORT MAP(module2_48_todown, module2_49_fromdown, clock, hardcoded_49, module2_48_fromdown, module2_49_todown); 
module2op_50: module2 PORT MAP(module2_49_todown, module2_50_fromdown, clock, hardcoded_50, module2_49_fromdown, module2_50_todown); 
module2op_51: module2 PORT MAP(module2_50_todown, module2_51_fromdown, clock, hardcoded_51, module2_50_fromdown, module2_51_todown); 
module2op_52: module2 PORT MAP(module2_51_todown, module2_52_fromdown, clock, hardcoded_52, module2_51_fromdown, module2_52_todown); 
module2op_53: module2 PORT MAP(module2_52_todown, module2_53_fromdown, clock, hardcoded_53, module2_52_fromdown, module2_53_todown); 
module2op_54: module2 PORT MAP(module2_53_todown, module2_54_fromdown, clock, hardcoded_54, module2_53_fromdown, module2_54_todown); 
module2op_55: module2 PORT MAP(module2_54_todown, module2_55_fromdown, clock, hardcoded_55, module2_54_fromdown, module2_55_todown); 
module2op_56: module2 PORT MAP(module2_55_todown, module2_56_fromdown, clock, hardcoded_56, module2_55_fromdown, module2_56_todown); 
module2op_57: module2 PORT MAP(module2_56_todown, module2_57_fromdown, clock, hardcoded_57, module2_56_fromdown, module2_57_todown); 
module2op_58: module2 PORT MAP(module2_57_todown, module2_58_fromdown, clock, hardcoded_58, module2_57_fromdown, module2_58_todown); 
module2op_59: module2 PORT MAP(module2_58_todown, module2_59_fromdown, clock, hardcoded_59, module2_58_fromdown, module2_59_todown); 
module2op_60: module2 PORT MAP(module2_59_todown, module2_60_fromdown, clock, hardcoded_60, module2_59_fromdown, module2_60_todown); 
module2op_61: module2 PORT MAP(module2_60_todown, module2_61_fromdown, clock, hardcoded_61, module2_60_fromdown, module2_61_todown); 
module2op_62: module2 PORT MAP(module2_61_todown, module2_62_fromdown, clock, hardcoded_62, module2_61_fromdown, module2_62_todown); 
module2op_63: module2 PORT MAP(module2_62_todown, module2_63_fromdown, clock, hardcoded_63, module2_62_fromdown, module2_63_todown); 
module2op_64: module2 PORT MAP(module2_63_todown, module2_64_fromdown, clock, hardcoded_64, module2_63_fromdown, module2_64_todown); 
module2op_65: module2 PORT MAP(module2_64_todown, module2_65_fromdown, clock, hardcoded_65, module2_64_fromdown, module2_65_todown); 
module2op_66: module2 PORT MAP(module2_65_todown, module2_66_fromdown, clock, hardcoded_66, module2_65_fromdown, module2_66_todown); 
module2op_67: module2 PORT MAP(module2_66_todown, module2_67_fromdown, clock, hardcoded_67, module2_66_fromdown, module2_67_todown); 
module2op_68: module2 PORT MAP(module2_67_todown, module2_68_fromdown, clock, hardcoded_68, module2_67_fromdown, module2_68_todown); 
module2op_69: module2 PORT MAP(module2_68_todown, module2_69_fromdown, clock, hardcoded_69, module2_68_fromdown, module2_69_todown); 
module2op_70: module2 PORT MAP(module2_69_todown, module2_70_fromdown, clock, hardcoded_70, module2_69_fromdown, module2_70_todown); 
module2op_71: module2 PORT MAP(module2_70_todown, module2_71_fromdown, clock, hardcoded_71, module2_70_fromdown, module2_71_todown); 
module2op_72: module2 PORT MAP(module2_71_todown, module2_72_fromdown, clock, hardcoded_72, module2_71_fromdown, module2_72_todown); 
module2op_73: module2 PORT MAP(module2_72_todown, module2_73_fromdown, clock, hardcoded_73, module2_72_fromdown, module2_73_todown); 
module2op_74: module2 PORT MAP(module2_73_todown, module2_74_fromdown, clock, hardcoded_74, module2_73_fromdown, module2_74_todown); 
module2op_75: module2 PORT MAP(module2_74_todown, module2_75_fromdown, clock, hardcoded_75, module2_74_fromdown, module2_75_todown); 
module2op_76: module2 PORT MAP(module2_75_todown, module2_76_fromdown, clock, hardcoded_76, module2_75_fromdown, module2_76_todown); 
module2op_77: module2 PORT MAP(module2_76_todown, module2_77_fromdown, clock, hardcoded_77, module2_76_fromdown, module2_77_todown); 
module2op_78: module2 PORT MAP(module2_77_todown, module2_78_fromdown, clock, hardcoded_78, module2_77_fromdown, module2_78_todown); 
module2op_79: module2 PORT MAP(module2_78_todown, module2_79_fromdown, clock, hardcoded_79, module2_78_fromdown, module2_79_todown); 
module2op_80: module2 PORT MAP(module2_79_todown, module2_80_fromdown, clock, hardcoded_80, module2_79_fromdown, module2_80_todown); 
module2op_81: module2 PORT MAP(module2_80_todown, module2_81_fromdown, clock, hardcoded_81, module2_80_fromdown, module2_81_todown); 
module2op_82: module2 PORT MAP(module2_81_todown, module2_82_fromdown, clock, hardcoded_82, module2_81_fromdown, module2_82_todown); 
module2op_83: module2 PORT MAP(module2_82_todown, module2_83_fromdown, clock, hardcoded_83, module2_82_fromdown, module2_83_todown); 
module2op_84: module2 PORT MAP(module2_83_todown, module2_84_fromdown, clock, hardcoded_84, module2_83_fromdown, module2_84_todown); 
module2op_85: module2 PORT MAP(module2_84_todown, module2_85_fromdown, clock, hardcoded_85, module2_84_fromdown, module2_85_todown); 
module2op_86: module2 PORT MAP(module2_85_todown, module2_86_fromdown, clock, hardcoded_86, module2_85_fromdown, module2_86_todown); 
module2op_87: module2 PORT MAP(module2_86_todown, module2_87_fromdown, clock, hardcoded_87, module2_86_fromdown, module2_87_todown); 
module2op_88: module2 PORT MAP(module2_87_todown, module2_88_fromdown, clock, hardcoded_88, module2_87_fromdown, module2_88_todown); 
module2op_89: module2 PORT MAP(module2_88_todown, module2_89_fromdown, clock, hardcoded_89, module2_88_fromdown, module2_89_todown); 
module2op_90: module2 PORT MAP(module2_89_todown, module2_90_fromdown, clock, hardcoded_90, module2_89_fromdown, module2_90_todown); 
module2op_91: module2 PORT MAP(module2_90_todown, module2_91_fromdown, clock, hardcoded_91, module2_90_fromdown, module2_91_todown); 
module2op_92: module2 PORT MAP(module2_91_todown, module2_92_fromdown, clock, hardcoded_92, module2_91_fromdown, module2_92_todown); 
module2op_93: module2 PORT MAP(module2_92_todown, module2_93_fromdown, clock, hardcoded_93, module2_92_fromdown, module2_93_todown); 
module2op_94: module2 PORT MAP(module2_93_todown, module2_94_fromdown, clock, hardcoded_94, module2_93_fromdown, module2_94_todown); 
module2op_95: module2 PORT MAP(module2_94_todown, module2_95_fromdown, clock, hardcoded_95, module2_94_fromdown, module2_95_todown); 
module2op_96: module2 PORT MAP(module2_95_todown, module2_96_fromdown, clock, hardcoded_96, module2_95_fromdown, module2_96_todown); 
module2op_97: module2 PORT MAP(module2_96_todown, module2_97_fromdown, clock, hardcoded_97, module2_96_fromdown, module2_97_todown); 
module2op_98: module2 PORT MAP(module2_97_todown, module2_98_fromdown, clock, hardcoded_98, module2_97_fromdown, module2_98_todown); 
module2op_99: module2 PORT MAP(module2_98_todown, module2_99_fromdown, clock, hardcoded_99, module2_98_fromdown, module2_99_todown); 
module2op_100: module2 PORT MAP(module2_99_todown, module2_100_fromdown, clock, hardcoded_100, module2_99_fromdown, module2_100_todown); 
module2op_101: module2 PORT MAP(module2_100_todown, module2_101_fromdown, clock, hardcoded_101, module2_100_fromdown, module2_101_todown); 
module2op_102: module2 PORT MAP(module2_101_todown, module2_102_fromdown, clock, hardcoded_102, module2_101_fromdown, module2_102_todown); 
module2op_103: module2 PORT MAP(module2_102_todown, module2_103_fromdown, clock, hardcoded_103, module2_102_fromdown, module2_103_todown); 
module2op_104: module2 PORT MAP(module2_103_todown, module2_104_fromdown, clock, hardcoded_104, module2_103_fromdown, module2_104_todown); 
module2op_105: module2 PORT MAP(module2_104_todown, module2_105_fromdown, clock, hardcoded_105, module2_104_fromdown, module2_105_todown); 
module2op_106: module2 PORT MAP(module2_105_todown, module2_106_fromdown, clock, hardcoded_106, module2_105_fromdown, module2_106_todown); 
module2op_107: module2 PORT MAP(module2_106_todown, module2_107_fromdown, clock, hardcoded_107, module2_106_fromdown, module2_107_todown); 
module2op_108: module2 PORT MAP(module2_107_todown, module2_108_fromdown, clock, hardcoded_108, module2_107_fromdown, module2_108_todown); 
module2op_109: module2 PORT MAP(module2_108_todown, module2_109_fromdown, clock, hardcoded_109, module2_108_fromdown, module2_109_todown); 
module2op_110: module2 PORT MAP(module2_109_todown, module2_110_fromdown, clock, hardcoded_110, module2_109_fromdown, module2_110_todown); 
module2op_111: module2 PORT MAP(module2_110_todown, module2_111_fromdown, clock, hardcoded_111, module2_110_fromdown, module2_111_todown); 
module2op_112: module2 PORT MAP(module2_111_todown, module2_112_fromdown, clock, hardcoded_112, module2_111_fromdown, module2_112_todown); 
module2op_113: module2 PORT MAP(module2_112_todown, module2_113_fromdown, clock, hardcoded_113, module2_112_fromdown, module2_113_todown); 
module2op_114: module2 PORT MAP(module2_113_todown, module2_114_fromdown, clock, hardcoded_114, module2_113_fromdown, module2_114_todown); 
module2op_115: module2 PORT MAP(module2_114_todown, module2_115_fromdown, clock, hardcoded_115, module2_114_fromdown, module2_115_todown); 
module2op_116: module2 PORT MAP(module2_115_todown, module2_116_fromdown, clock, hardcoded_116, module2_115_fromdown, module2_116_todown); 
module2op_117: module2 PORT MAP(module2_116_todown, module2_117_fromdown, clock, hardcoded_117, module2_116_fromdown, module2_117_todown); 
module2op_118: module2 PORT MAP(module2_117_todown, module2_118_fromdown, clock, hardcoded_118, module2_117_fromdown, module2_118_todown); 
module2op_119: module2 PORT MAP(module2_118_todown, module2_119_fromdown, clock, hardcoded_119, module2_118_fromdown, module2_119_todown); 
module2op_120: module2 PORT MAP(module2_119_todown, module2_120_fromdown, clock, hardcoded_120, module2_119_fromdown, module2_120_todown); 
module2op_121: module2 PORT MAP(module2_120_todown, module2_121_fromdown, clock, hardcoded_121, module2_120_fromdown, module2_121_todown); 
module2op_122: module2 PORT MAP(module2_121_todown, module2_122_fromdown, clock, hardcoded_122, module2_121_fromdown, module2_122_todown); 
module2op_123: module2 PORT MAP(module2_122_todown, module2_123_fromdown, clock, hardcoded_123, module2_122_fromdown, module2_123_todown); 
module2op_124: module2 PORT MAP(module2_123_todown, module2_124_fromdown, clock, hardcoded_124, module2_123_fromdown, module2_124_todown); 
module2op_125: module2 PORT MAP(module2_124_todown, module2_125_fromdown, clock, hardcoded_125, module2_124_fromdown, module2_125_todown); 
module2op_126: module2 PORT MAP(module2_125_todown, module2_126_fromdown, clock, hardcoded_126, module2_125_fromdown, module2_126_todown); 
module3op: module3 PORT MAP(module2_126_todown, clock, hardcoded_127, module2_126_fromdown); 
end Behavioral; 

