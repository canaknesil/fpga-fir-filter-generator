VHDL code has hot been implemented yet.
Filter signal: [ 5 ]

